
DATAPATH
-- Author: Nguyễn Kiêm Hùng
LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
use work.User_Lib.all;
use ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
--use ieee.numeric_std.all;
ENTITY Datapath IS
   GENERIC (
            DATA_WIDTH        :     integer   := 8;     -- Word Width
            ADDR_WIDTH        :     integer   := 2      -- Address width
           
    );
   PORT ( Clock, Reset: IN STD_LOGIC ;
          Start: IN STD_LOGIC ;
          
          Min_Sel, Addr_Sel: IN STD_LOGIC; -- The signal selects the input data and address for memory
          Int_WE, WE: IN STD_LOGIC;
          Int_RE, RE: IN STD_LOGIC;
          
          LD_i, LD_j: IN STD_LOGIC; -- Load signal for Counter i
          En_i, En_j: IN STD_LOGIC;
          EN_A, EN_B: IN STD_LOGIC;
          data_in : IN STD_LOGIC_VECTOR (DATA_WIDTH - 1 downto 0);
          addr_in : IN STD_LOGIC_VECTOR (ADDR_WIDTH - 1 downto 0);
          Zi,Zj : OUT STD_LOGIC;
	        A_gt_B : OUT STD_LOGIC;
	        data_out : OUT STD_LOGIC_VECTOR (DATA_WIDTH - 1 downto 0) ) ;
   END Datapath ;

ARCHITECTURE RTL OF Datapath IS
  CONSTANT K   : integer   := 2**ADDR_WIDTH;
  --TYPE State_type IS (A, B, C) ;
  SIGNAL State : STD_LOGIC_VECTOR(4 DOWNTO 0) ;
  -- Signal for connecting to Mem_block
  signal nReset :      std_logic := '0';
  signal addr : std_logic_vector( ADDR_WIDTH-1 downto 0);
  signal  wen  :       std_logic;
  signal  datain :  std_logic_vector(DATA_WIDTH -1 downto 0);
  signal  ren :       std_logic;
  signal i,i_plus_1,j,i_mux_j : std_logic_vector( ADDR_WIDTH-1 downto 0);
  signal A,B,A_mux_B : std_logic_vector(DATA_WIDTH -1 downto 0);
  signal dataout :   std_logic_vector(DATA_WIDTH -1 downto 0);
BEGIN
  nReset <= not Reset;
  i_mux_j <= i when addr_sel = '0' else j;
  A_mux_B <= A when Min_sel = '0' else B;
  addr <= ADDR_in when Start = '0' else i_mux_j;
  datain <= data_in when Start = '0' else A_mux_B;
  wen <= int_WE or WE;
  ren <= int_RE or RE;
 -- Memory block
 Mem_Block:  dpmem
    generic map
    (
      DATA_WIDTH => DATA_WIDTH,
      ADDR_WIDTH => ADDR_WIDTH
      )
     
     port map (
       
      clk      => clock,
      nReset   => nReset,
      addr     => addr,
      Wen      => wen,
      Datain   => datain,
      
      Ren      => ren,
      
      Dataout  => dataout
      
      );
  --------------
  -- Register A
  RegA: regn
  generic map
     (
      N => DATA_WIDTH
      )
    port map (
      D => dataout, 
      Reset   => Reset,
      clock   => clock,
      En      => En_A,
      Q  => A
      
      );  
  -- Register B
  RegB: regn
  generic map
     (
      N => DATA_WIDTH
      )
    port map (
      D => dataout, 
      Reset   => Reset,
      clock   => clock,
      En      => En_B,
      Q  => B
      
      );     
 -- Comrator A>B
 A_gt_B <= '1' WHEN A>B ELSE '0';     
-- Counter i
Cnt_i: Counter_n
  generic map
     (
      N => ADDR_WIDTH
      )
    port map (
      clk   => clock,
      Reset   => Reset,
      Enable  => En_i,
      Load    => LD_i,
      Din => (OTHERS => '0'), 
      Count  => i
       ); 
  zi <= '0' WHEN i < conv_std_logic_vector(K-1,ADDR_WIDTH) ELSE '1';      
-- Counter j
Cnt_j: Counter_n
  generic map
     (
      N => ADDR_WIDTH
      )
    port map (
      clk   => clock,
      Reset   => Reset,
      Enable  => En_j,
      Load    => LD_j,
      Din => i_plus_1, 
      Count  => j
       ); 
  i_plus_1 <= i + 1;
  zj <= '0' WHEN j /= conv_std_logic_vector(0,ADDR_WIDTH) ELSE '1';      
  -- Output
    data_out <= Dataout;
    
END RTL;   

LIB USER
--This confidential and proprietary software may be used
--only as authorized by a licensing agreement from
--Laboratory for Smart Integrated Systems (SIS), VNU University of Engineering and Technology (VNU-UET).
-- (C) COPYRIGHT 2015
-- ALL RIGHTS RESERVED
-- The entire notice above must be reproduced on all authorized copies.
--
-- Filename : RCA_define.v
-- Author : Hung Nguyen
-- Date : 
-- Version : 0.1
-- Description Package declares all constants, types, 
-- and components for project.               
-- Modification History:
-- Date By Version Change Description
-- ========================================================
-- 05/08.2014  0.1 Original
-- ========================================================
library IEEE;
use IEEE.std_logic_1164.all;
USE ieee.numeric_std.all ;
use std.textio.all;

package User_Lib is

-- Constant for datapath
  Constant   DATA_WIDTH  :     integer   := 16;     -- Word Width
  Constant   ADDR_WIDTH  :     integer   := 16 ;     -- Address width
--constant PORT_NUM : integer := 5;

-- Type Definition
   -- type ADDR_ARRAY_TYPE is array (VC_NUM-1 DOWNTO 0) of std_logic_vector (ADDR_WIDTH-1 downto 0);
   

-- **************************************************************
--COMPONENTs
--------------------------------
-- FULL ADDER 1 bit
COMPONENT fulladder_1b 

    PORT (
        x,y :  IN  std_logic;
        cin :  IN  std_logic;
        s   :  OUT std_logic;
        cout : OUT std_logic);
END COMPONENT;

-------------------------------------------
component dpmem 
   generic (
     DATA_WIDTH        :     integer   := 16;     -- Word Width
     ADDR_WIDTH        :     integer   := 16      -- Address width
     );
 
   port (
     -- Writing
     Clk              : in  std_logic;          -- clock
     nReset             : in  std_logic; -- Reset input
     addr              : in  std_logic_vector(ADDR_WIDTH -1 downto 0);   --  Address
     -- Writing Port
     Wen               : in  std_logic;          -- Write Enable
     Datain            : in  std_logic_vector(DATA_WIDTH -1 downto 0) := (others => '0');   -- Input Data
     -- Reading Port
     
     Ren               : in  std_logic;          -- Read Enable
     Dataout           : out std_logic_vector(DATA_WIDTH -1 downto 0)   -- Output data
     
     );
  
  end component;
--------------------------------------------  
COMPONENT regn 
  GENERIC (N : INTEGER := 16);
  PORT (
      D : IN STD_LOGIC_VECTOR (N-1 DOWNTO 0) ;
   	  Reset, Clock, En : IN STD_LOGIC ;
	    Q : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	    );
END COMPONENT ;
----------------------------------------------
COMPONENT counter_n 
    GENERIC (N : Integer := 2);
		PORT (clk:  IN std_logic;
			  reset: IN std_logic;
			  enable: IN std_logic;
			  Load : IN std_logic;
			  Din  : IN std_logic_vector(N-1 downto 0);
			  count:  OUT std_logic_vector(N-1 downto 0));
END COMPONENT;
--------------------------------------------------
COMPONENT Sorter 
   GENERIC (
            DATA_WIDTH        :     integer   := 8;     -- Word Width
            ADDR_WIDTH        :     integer   := 2      -- Address width
           
    );
   PORT ( Clock, nReset: IN STD_LOGIC ;
          Start: IN STD_LOGIC ;
          
          WE: IN STD_LOGIC;
          RE: IN STD_LOGIC;
          
          data_in : IN STD_LOGIC_VECTOR (DATA_WIDTH - 1 downto 0);
          addr_in : IN STD_LOGIC_VECTOR (ADDR_WIDTH - 1 downto 0);
          Done    : OUT STD_LOGIC;
	        data_out : OUT STD_LOGIC_VECTOR (DATA_WIDTH - 1 downto 0) ) ;
   END COMPONENT ;
---------------------------------------------------
COMPONENT Controller 
   PORT ( Clock, nReset: IN STD_LOGIC ;
          Start: IN STD_LOGIC ;
          
          Zi, Zj: IN STD_LOGIC; -- Output signal of Comparator i
          A_gt_B: IN STD_LOGIC;
          
          Addr_sel, Min_sel, int_RE, int_WE: OUT STD_LOGIC; 
          LD_i, LD_j: OUT STD_LOGIC; -- Load signal for Counter i
          En_i, En_j: OUT STD_LOGIC;
          EN_A, EN_B: OUT STD_LOGIC;
          reset : OUT STD_LOGIC;
	        Done : OUT STD_LOGIC ) ;
   END COMPONENT ;
----------------------------------
COMPONENT Datapath 
   GENERIC (
            DATA_WIDTH        :     integer   := 8;     -- Word Width
            ADDR_WIDTH        :     integer   := 2      -- Address width
           
    );
   PORT ( Clock, Reset: IN STD_LOGIC ;
          Start: IN STD_LOGIC ;
          
          Min_Sel, Addr_Sel: IN STD_LOGIC; -- The signal selects the input data and address for memory
          Int_WE, WE: IN STD_LOGIC;
          Int_RE, RE: IN STD_LOGIC;
          
          LD_i, LD_j: IN STD_LOGIC; -- Load signal for Counter i
          En_i, En_j: IN STD_LOGIC;
          EN_A, EN_B: IN STD_LOGIC;
          data_in : IN STD_LOGIC_VECTOR (DATA_WIDTH - 1 downto 0);
          addr_in : IN STD_LOGIC_VECTOR (ADDR_WIDTH - 1 downto 0);
          Zi,Zj : OUT STD_LOGIC;
	        A_gt_B : OUT STD_LOGIC;
	        data_out : OUT STD_LOGIC_VECTOR (DATA_WIDTH - 1 downto 0) ) ;
   END COMPONENT;
-----------------------------------------
COMPONENT xor2 
  PORT(
       I1   : IN STD_LOGIC;
       I2   : IN STD_LOGIC;
       Y   : OUT STD_LOGIC);
END COMPONENT;

------------------------------------------------------
Component mux4to1 
   Generic ( 
		    DATA_WIDTH : integer := 8);
   PORT (A, B, C, D: IN  	std_logic_vector (DATA_WIDTH-1 downto 0);
        SEL : IN 	 std_logic_vector (1 downto 0);
        Z: OUT 	std_logic_vector (DATA_WIDTH-1 downto 0)
               );
END Component;
-----------------
-- You need to add the other components here......
-----------------
end User_Lib;

PACKAGE BODY User_Lib IS
	-- package body declarations

END PACKAGE BODY User_Lib;

DPMEM
-- Author: Nguyễn Kiêm Hùng
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
 
-------------------------------------------------------------------------------
-- Synchronous Dual Port Memory
-------------------------------------------------------------------------------
entity dpmem is
  generic (
    DATA_WIDTH        :     integer   := 16;     -- Word Width
    ADDR_WIDTH        :     integer   := 16      -- Address width
    );

  port (
    -- Writing
    Clk              : in  std_logic;          -- clock
	nReset             : in  std_logic; -- Reset input
    addr              : in  std_logic_vector(ADDR_WIDTH -1 downto 0);   --  Address
	-- Writing Port
	Wen               : in  std_logic;          -- Write Enable
    Datain            : in  std_logic_vector(DATA_WIDTH -1 downto 0) := (others => '0');   -- Input Data
    -- Reading Port
    
    Ren               : in  std_logic;          -- Read Enable
    Dataout           : buffer std_logic_vector(DATA_WIDTH -1 downto 0)   -- Output data
    
    );
end dpmem;
 
architecture dpmem_arch of dpmem is
   
  type DATA_ARRAY is array (integer range <>) of std_logic_vector(DATA_WIDTH -1 downto 0); -- Memory Type
  signal   M       :     DATA_ARRAY(0 to (2**ADDR_WIDTH) -1) := (others => (others => '0'));  -- Memory model
-- you can add more code for your application by increase the PM_Size

begin  -- dpmem_arch
	
	
  --  Read/Write process

  RW_Proc : process (clk, nReset)
  begin  
    if nReset = '0' then
          Dataout <= (others => '0');
          M <= (others => (others => '0')); -- initialize memory
    elsif (clk'event and clk = '1') then   -- rising clock edge
        if Wen = '1' then
			   M(conv_integer(addr))      <= Datain; -- ensure that data cant overwrite on program
        else
			   if Ren = '1' then
				    Dataout <= M(conv_integer(addr));
			   else
				   Dataout <= Dataout;
			   end if;
		   end if;
      end if;
  end process  RW_Proc;
     
end dpmem_arch;

REGn
-- Author: Nguyễn Kiêm Hùng
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.User_Lib.all;
ENTITY regn IS
  GENERIC (N : INTEGER := 16);
  PORT (
      D : IN STD_LOGIC_VECTOR (N-1 DOWNTO 0) ;
   	  Reset, Clock, En : IN STD_LOGIC ;
	    Q : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	    );
END regn ;
ARCHITECTURE Behavior OF regn IS
  BEGIN
    PROCESS (Reset, Clock)
      BEGIN
        IF RESET='1' THEN
          Q <= (OTHERS => '0');
        ELSIF (CLOCK'EVENT AND CLOCK='1') THEN
          IF (EN = '1') THEN
            Q <= D;
          END IF;
        END IF;

   END PROCESS ;
END Behavior ;

COUNTER
-- Author: Nguyễn Kiêm Hùng
--counter.vhd
library ieee ;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
ENTITY counter_n IS 
    GENERIC (N : Integer := 2);
		PORT (clk:  IN std_logic;
			  reset: IN std_logic;
			  enable: IN std_logic;
			  Load : IN std_logic;
			  Din  : IN std_logic_vector(N-1 downto 0);
			  count:  OUT std_logic_vector(N-1 downto 0));
END counter_n;
ARCHITECTURE behav OF counter_n IS
  SIGNAL pre_count: std_logic_vector(N-1 downto 0);  BEGIN
    PROCESS(clk, enable, reset)
		    BEGIN
		      IF reset = '1' THEN
		        pre_count <= (OTHERS =>'0');
		      ELSIF (clk='1' and clk'event) THEN
		        IF Load = '1' THEN
		            pre_count <= Din;
		        ELSIF enable = '1' THEN
			          pre_count <= pre_count + "1"; 
			          
			       END IF;
		 	  END IF;
    END PROCESS;
    count <= pre_count;
END behav;

CONTROLER
-- Author: Nguyễn Kiêm Hùng
LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
use work.User_Lib.all;
ENTITY Controller IS
   PORT ( Clock, nReset: IN STD_LOGIC ;
          Start: IN STD_LOGIC ;
          
          Zi, Zj: IN STD_LOGIC; -- Output signal of Comparator i
          A_gt_B: IN STD_LOGIC;
          
          Addr_sel, Min_sel, int_RE, int_WE: OUT STD_LOGIC; 
          LD_i, LD_j: OUT STD_LOGIC; -- Load signal for Counter i
          En_i, En_j: OUT STD_LOGIC;
          EN_A, EN_B: OUT STD_LOGIC;
          reset : OUT STD_LOGIC;
	        Done : OUT STD_LOGIC ) ;
   END Controller ;
ARCHITECTURE Behavior OF Controller IS
  --TYPE State_type IS (A, B, C) ;
  SIGNAL State : STD_LOGIC_VECTOR(4 DOWNTO 0) ;
  SIGNAL EN_A_T: STD_LOGIC;
BEGIN
-- State transitions 
  PROCESS ( nReset, Clock )
    BEGIN
      
      IF nReset = '0' THEN
	       STATE <= "00000" ; -- STATE 0
      ELSIF (Clock'EVENT AND Clock = '1') THEN
        CASE STATE IS
           WHEN "00000" =>
               STATE <= "00001"; -- STATE 1
           WHEN "00001" =>    
               IF START = '1' THEN
	               STATE <= "00010"; -- STATE 2
	             ELSE
	               STATE <= "00001"; -- STATE 1
               END IF ;
            WHEN "00010" =>
                STATE <= "00011"; -- STATE 3
            WHEN "00011" =>
                IF Zi = '0' THEN
                  STATE <= "00100"; -- STATE 4
                ELSE
                  STATE <= "10001"; -- STATE 17
                END IF ;
             WHEN "00100" => --4
                STATE <= "00110"; -- STATE 5
             WHEN "00101" => --5
                STATE <= "00110"; -- STATE 6
             WHEN "00110" => --6
                STATE <= "00111"; -- STATE 7   
             WHEN "00111" =>
                IF Zj = '0' THEN
                  STATE <= "01000"; -- STATE 8
                ELSE
                  STATE <= "10000"; -- STATE 16
                END IF ;  
             WHEN "01000" =>  --8  
                STATE <= "01001"; -- STATE 9 
             WHEN "01001" => --9
                STATE <= "01010"; -- STATE 10 
             WHEN "01010" => --10   
                IF A_gt_B = '1' THEN
                  STATE <= "01011"; -- STATE 11
                ELSE
                  STATE <= "01111"; -- STATE 15
                END IF ; 
             WHEN "01011" => 
                STATE <= "01100"; -- STATE 12
             WHEN "01100" => 
                STATE <= "01101"; -- STATE 13
             WHEN "01101" => -- 13
                STATE <= "01111"; -- STATE 14
             WHEN "01110" => --14
                STATE <= "01111"; -- STATE 15
             WHEN "01111" => --15
                STATE <= "00111"; -- STATE 7
             WHEN "10000" => 
                STATE <= "00011"; -- STATE 3  
             WHEN "10001" => 
                STATE <= "10010"; -- STATE 18 
             WHEN "10010" => 
                STATE <= "10011"; -- STATE 3                              
            WHEN OTHERs =>
                STATE <= "00001"; -- STATE 1 
          END CASE ;
  END IF ;


  END PROCESS ;
-- Output function
  -- Clear Registers
   Reset <= '1' WHEN STATE = "00000" ELSE '0' ;
  -- Load data into counters  
   LD_i <= '1' WHEN STATE = "00010" ELSE '0' ;
   LD_j <= '1' WHEN STATE = "00110" ELSE '0' ;
 -- Enable Counters
   EN_i <= '1' WHEN STATE = "10000" ELSE '0' ;
   EN_j <= '1' WHEN STATE = "01111" ELSE '0' ;  
 WITH STATE SELECT   
	 	Addr_sel <= '0' when "00100"|"01011"|"01101",
		    	       '1' when "01000"|"01100",
		    	
		    	       '0' when OTHERS;
  WITH STATE SELECT   
	 	Min_sel <= '0' when "01100",
		    	      '1' when "01011",
		    	
		    	       '0' when OTHERS;		    	       
 WITH STATE SELECT   
	 	Int_RE <= '1' when "00100"|"01000"|"01101",
		    	        	
		    	     '0' when OTHERS;
 WITH STATE SELECT   
	 	Int_WE <= '1' when "01011"|"01100",
		    	        	
		    	     '0' when OTHERS;	
 WITH STATE SELECT   
	 	EN_A_T <= '1' when "00100"|"01101",
		    	        	
		    	     '0' when OTHERS;		
EN_A_PRoC: PROCESS ( nReset, Clock )
    BEGIN 
      IF nReset = '0' THEN
	       EN_A <= '0' ; 
      ELSIF (Clock'EVENT AND Clock = '1') THEN
         EN_A <= EN_A_T;
    END IF;
END PROCESS ;       
 EN_B <= '1' WHEN STATE = "01001" ELSE '0' ;		 
 Done <= '1' WHEN (STATE = "10001") OR (STATE = "10010") ELSE '0' ;		    	     	    	     	    	     
END Behavior;   

SORTER
-- Author: Nguyễn Kiêm Hùng
LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
use work.User_Lib.all;
USE ieee.std_logic_unsigned.all;

ENTITY Sorter IS
   GENERIC (
            DATA_WIDTH        :     integer   := 8;     -- Word Width
            ADDR_WIDTH        :     integer   := 2      -- Address width
           
    );
   PORT ( Clock, nReset: IN STD_LOGIC ;
          Start: IN STD_LOGIC ;
          
          WE: IN STD_LOGIC;
          RE: IN STD_LOGIC;
          
          data_in : IN STD_LOGIC_VECTOR (DATA_WIDTH - 1 downto 0);
          addr_in : IN STD_LOGIC_VECTOR (ADDR_WIDTH - 1 downto 0);
          Done    : OUT STD_LOGIC;
	        data_out : OUT STD_LOGIC_VECTOR (DATA_WIDTH - 1 downto 0) ) ;
   END Sorter ;
ARCHITECTURE RTL OF Sorter IS
  SIGNAL Min_Sel, Addr_Sel: STD_LOGIC;
  SIGNAL  Int_RE, Int_WE: STD_LOGIC;
  SIGNAL LD_i, LD_j:  STD_LOGIC; -- Load signal for Counter i
  SIGNAL En_i, En_j:  STD_LOGIC;
  SIGNAL EN_A, EN_B:  STD_LOGIC; 
  SIGNAL Zi,Zj : STD_LOGIC;  
  SIGNAL A_gt_B : STD_LOGIC;
	SIGNAL Reset : STD_LOGIC;     
BEGIN
CRTL_U: Controller 
   PORT MAP( Clock,
             nReset,
             Start,
          
          Zi,
          Zj, -- Output signal of Comparator i
          A_gt_B,
          
          Addr_sel,
          Min_sel,
          int_RE,
          int_WE, 
          LD_i,
          LD_j, -- Load signal for Counter i
          En_i,
          En_j,
          EN_A,
          EN_B,
          reset,
	        Done) ;
   
Datapath_U: Datapath
  GENERIC MAP(
            DATA_WIDTH => DATA_WIDTH,     -- Word Width
            ADDR_WIDTH => ADDR_WIDTH      -- Address width
           
          )
   PORT MAP( Clock, 
          Reset,
          Start,
          
          Min_Sel, 
          Addr_Sel, -- The signal selects the input data and address for memory
          Int_WE, 
          WE,
          Int_RE, 
          RE,
          
          LD_i, 
          LD_j, -- Load signal for Counter i
          En_i,
          En_j,
          EN_A,
          EN_B,
          data_in,
          addr_in,
          Zi,
          Zj,
	        A_gt_B,
	        data_out ) ;
END RTL;  